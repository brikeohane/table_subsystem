library ieee;
use ieee.std_logic_1164.all; 

entity read_fsm is
	port(
		clk, reset: in std_logic;
		start: 		in std_logic;
		key_in:		in std_logic_vector(47 downto 0);
		key_out:	out std_logic_vector(47 downto 0);
		data_in: 	in std_logic_vector(1 downto 0);
		hit_in:		in std_logic;
		data_out:	out std_logic_vector(1 downto 0);
		hit_out:	out std_logic;
		done:		out std_logic
	);
end read_fsm;

architecture read_fsm_rtl of read_fsm is

	type state_type is (initial, reading, finished);
	signal state_reg, state_next: state_type;
	signal key_reg: std_logic_vector(47 downto 0);
	signal data_reg: std_logic_vector(1 downto 0);
	signal hit_reg: std_logic;

begin

	-- Update the current state every clock cycle
	STATE_REGISTER: process(clk,reset) 
	begin
		if(reset = '1') then 
			state_reg <= initial;
		elsif (clk'event and clk = '1') then 
			state_reg <= state_next;
		end if;
	end process;

	INPUT_REGISTER: process(clk,key_in,data_in)
	begin
		if(clk'event and clk = '1') then 
			key_reg <= key_in;
			data_reg <= data_in;
			hit_reg <= hit_in;
		end if;
	end process;

	-- Define state transitions for the FSM
	NEXT_STATE: process(state_reg, start) 
	begin
		case state_reg is 
			when initial =>
				if (start = '1') then 
					state_next <= reading;
				else
					state_next <= initial;
				end if; 
			when reading =>
				state_next <= finished;
			when finished => 
				state_next <= initial;
		end case;
	end process;

	-- Specify Moore outputs for the FSM
	STATE_OUTPUT: process(state_reg)
	begin
		if(state_reg = finished) then
			done <= '1';
		else
			done <= '0'; 
		end if;
	end process;

	-- Output to CAM
	key_out <= key_reg;

	-- Output to Interface
	data_out <= data_reg;
	hit_out <= hit_reg;
end read_fsm_rtl;










